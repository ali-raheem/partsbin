/*
   Copyright 2020 Ali Raheem <github@shoryuken.me>

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and limitations under the License.
*/

module mux (a, b, q, switch);
   parameter BUS_WIDTH = 4;
   input [BUS_WIDTH - 1:0] a;
   input [BUS_WIDTH - 1:0] b;
   output [BUS_WIDTH - 1:0] q;
   input 		   switch;

   assign q = switch ? a : b;
   
endmodule // mux
