/*
   Copyright 2018 Ali Raheem <ali.raheem@gmail.com>

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and limitations under the License.
*/

module sseg_tb ();
   reg [3:0] in;
   wire [6:0] out;
   reg 	      oe;

   sseg DUT(
	    .in(in),
	    .out_q(out),
	    .oe(oe)
	    );
   initial begin
      $dumpfile("sseg.vcd");
      $dumpvars(0, sseg_tb);
      in = 0;
      oe = 1;
      #100
	$finish;
   end
   always #5 in = in + 1;
endmodule // sseg_tb

   
   
